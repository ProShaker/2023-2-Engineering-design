** Profile: "SCHEMATIC1-Task1"  [ c:\users\kimhyeongjun\documents\github\2023-2-engineering-design\pspice\first\231001_ex1_first-PSpiceFiles\SCHEMATIC1\Task1.sim ] 

** Creating circuit file "Task1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\KimHyeongJun\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 20 1Hz 10kHz
.STEP PARAM C_E LIST 50uF, 100uF, 150uF, 200uF 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
