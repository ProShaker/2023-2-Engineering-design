** Profile: "SCHEMATIC1-Task2"  [ C:\Users\KimHyeongJun\Documents\GitHub\2023-2-Engineering-design\PSPICE\First\231001_ex2-PSpiceFiles\SCHEMATIC1\Task2.sim ] 

** Creating circuit file "Task2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\KimHyeongJun\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 20 100Hz 100MegHz
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
